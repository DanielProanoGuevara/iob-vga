   // VGA
      input  [11:0] rgb,
      output v_sync,
      output h_sync,
      output [3:0] Red,
      output [3:0] Green,
      output [3:0] Blue,
      output [9:0] pixel_x,
      output [9:0] pixel_y,
